library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity cos625_24bit is
	port( address : IN INTEGER := 0;
		 cosx : OUT std_logic_vector (23 downto 0));
end cos625_24bit;

architecture cos625_24bit_ARCH of cos625_24bit is
	type cosromarray is array (0 to 624) of std_logic_vector (23 downto 0);
	constant cosxrom : cosromarray := (
X"7FFFFF",
X"7FFE58",
X"7FF960",
X"7FF119",
X"7FE582",
X"7FD69C",
X"7FC468",
X"7FAEE5",
X"7F9615",
X"7F79F7",
X"7F5A8E",
X"7F37D8",
X"7F11D8",
X"7EE88F",
X"7EBBFD",
X"7E8C23",
X"7E5904",
X"7E229F",
X"7DE8F7",
X"7DAC0E",
X"7D6BE3",
X"7D287B",
X"7CE1D5",
X"7C97F4",
X"7C4AD9",
X"7BFA88",
X"7BA701",
X"7B5048",
X"7AF65D",
X"7A9945",
X"7A3900",
X"79D592",
X"796EFC",
X"790543",
X"789868",
X"78286E",
X"77B558",
X"773F2A",
X"76C5E5",
X"76498E",
X"75CA28",
X"7547B5",
X"74C23A",
X"7439B9",
X"73AE36",
X"731FB6",
X"728E3A",
X"71F9C8",
X"716263",
X"70C810",
X"702AD1",
X"6F8AAB",
X"6EE7A2",
X"6E41BB",
X"6D98FA",
X"6CED63",
X"6C3EFA",
X"6B8DC4",
X"6AD9C6",
X"6A2304",
X"696984",
X"68AD49",
X"67EE58",
X"672CB8",
X"66686C",
X"65A17A",
X"64D7E6",
X"640BB7",
X"633CF1",
X"626B9A",
X"6197B7",
X"60C14D",
X"5FE863",
X"5F0CFE",
X"5E2F22",
X"5D4ED8",
X"5C6C23",
X"5B870A",
X"5A9F92",
X"59B5C3",
X"58C9A1",
X"57DB33",
X"56EA80",
X"55F78C",
X"550260",
X"540B00",
X"531174",
X"5215C1",
X"5117EF",
X"501803",
X"4F1606",
X"4E11FC",
X"4D0BED",
X"4C03E0",
X"4AF9DC",
X"49EDE7",
X"48E008",
X"47D046",
X"46BEA9",
X"45AB38",
X"4495F8",
X"437EF3",
X"42662F",
X"414BB2",
X"402F86",
X"3F11B0",
X"3DF239",
X"3CD127",
X"3BAE82",
X"3A8A52",
X"39649F",
X"383D6F",
X"3714CA",
X"35EAB9",
X"34BF43",
X"339270",
X"326447",
X"3134D0",
X"300413",
X"2ED218",
X"2D9EE7",
X"2C6A88",
X"2B3503",
X"29FE5F",
X"28C6A6",
X"278DDE",
X"265410",
X"251945",
X"23DD84",
X"22A0D5",
X"216341",
X"2024CF",
X"1EE589",
X"1DA576",
X"1C649F",
X"1B230C",
X"19E0C5",
X"189DD3",
X"175A3D",
X"16160D",
X"14D14B",
X"138BFF",
X"124631",
X"10FFEA",
X"0FB933",
X"0E7213",
X"0D2A94",
X"0BE2BE",
X"0A9A99",
X"09522E",
X"080985",
X"06C0A6",
X"05779B",
X"042E6C",
X"02E521",
X"019BC3",
X"00525A",
X"FF08F0",
X"FDBF8C",
X"FC7636",
X"FB2CF8",
X"F9E3DA",
X"F89AE4",
X"F75220",
X"F60995",
X"F4C14B",
X"F3794C",
X"F231A1",
X"F0EA50",
X"EFA364",
X"EE5CE4",
X"ED16D8",
X"EBD14A",
X"EA8C42",
X"E947C8",
X"E803E4",
X"E6C09F",
X"E57E01",
X"E43C13",
X"E2FADD",
X"E1BA67",
X"E07ABA",
X"DF3BDD",
X"DDFDD9",
X"DCC0B7",
X"DB847E",
X"DA4936",
X"D90EE9",
X"D7D59D",
X"D69D5B",
X"D5662C",
X"D43016",
X"D2FB23",
X"D1C75A",
X"D094C3",
X"CF6367",
X"CE334C",
X"CD047B",
X"CBD6FB",
X"CAAAD6",
X"C98011",
X"C856B5",
X"C72ECA",
X"C60858",
X"C4E365",
X"C3BFFA",
X"C29E1E",
X"C17DD8",
X"C05F30",
X"BF422E",
X"BE26D9",
X"BD0D38",
X"BBF552",
X"BADF2F",
X"B9CAD6",
X"B8B84D",
X"B7A79D",
X"B698CC",
X"B58BE1",
X"B480E4",
X"B377DA",
X"B270CB",
X"B16BBE",
X"B068BA",
X"AF67C4",
X"AE68E5",
X"AD6C21",
X"AC7181",
X"AB790A",
X"AA82C3",
X"A98EB2",
X"A89CDE",
X"A7AD4D",
X"A6C004",
X"A5D50B",
X"A4EC67",
X"A4061E",
X"A32236",
X"A240B5",
X"A161A2",
X"A08501",
X"9FAAD8",
X"9ED32D",
X"9DFE06",
X"9D2B69",
X"9C5B59",
X"9B8DDE",
X"9AC2FC",
X"99FAB9",
X"993519",
X"987222",
X"97B1D9",
X"96F443",
X"963964",
X"958143",
X"94CBE2",
X"941948",
X"936978",
X"92BC77",
X"92124A",
X"916AF6",
X"90C67D",
X"9024E6",
X"8F8633",
X"8EEA69",
X"8E518C",
X"8DBBA0",
X"8D28A9",
X"8C98AA",
X"8C0BA8",
X"8B81A6",
X"8AFAA8",
X"8A76B0",
X"89F5C3",
X"8977E4",
X"88FD16",
X"88855C",
X"8810BA",
X"879F32",
X"8730C7",
X"86C57C",
X"865D54",
X"85F852",
X"859678",
X"8537C9",
X"84DC47",
X"8483F5",
X"842ED5",
X"83DCE9",
X"838E32",
X"8342B5",
X"82FA71",
X"82B569",
X"8273A0",
X"823515",
X"81F9CC",
X"81C1C6",
X"818D04",
X"815B87",
X"812D51",
X"810263",
X"80DABE",
X"80B664",
X"809554",
X"807790",
X"805D19",
X"8045F0",
X"803214",
X"802187",
X"801449",
X"800A5A",
X"8003BA",
X"80006A",
X"80006A",
X"8003BA",
X"800A5A",
X"801449",
X"802187",
X"803214",
X"8045F0",
X"805D19",
X"807790",
X"809554",
X"80B664",
X"80DABE",
X"810263",
X"812D51",
X"815B87",
X"818D04",
X"81C1C6",
X"81F9CC",
X"823515",
X"8273A0",
X"82B569",
X"82FA71",
X"8342B5",
X"838E32",
X"83DCE9",
X"842ED5",
X"8483F5",
X"84DC47",
X"8537C9",
X"859678",
X"85F852",
X"865D54",
X"86C57C",
X"8730C7",
X"879F32",
X"8810BA",
X"88855C",
X"88FD16",
X"8977E4",
X"89F5C3",
X"8A76B0",
X"8AFAA8",
X"8B81A6",
X"8C0BA8",
X"8C98AA",
X"8D28A9",
X"8DBBA0",
X"8E518C",
X"8EEA69",
X"8F8633",
X"9024E6",
X"90C67D",
X"916AF6",
X"92124A",
X"92BC77",
X"936978",
X"941948",
X"94CBE2",
X"958143",
X"963964",
X"96F443",
X"97B1D9",
X"987222",
X"993519",
X"99FAB9",
X"9AC2FC",
X"9B8DDE",
X"9C5B59",
X"9D2B69",
X"9DFE06",
X"9ED32D",
X"9FAAD8",
X"A08501",
X"A161A2",
X"A240B5",
X"A32236",
X"A4061E",
X"A4EC67",
X"A5D50B",
X"A6C004",
X"A7AD4D",
X"A89CDE",
X"A98EB2",
X"AA82C3",
X"AB790A",
X"AC7181",
X"AD6C21",
X"AE68E5",
X"AF67C4",
X"B068BA",
X"B16BBE",
X"B270CB",
X"B377DA",
X"B480E4",
X"B58BE1",
X"B698CC",
X"B7A79D",
X"B8B84D",
X"B9CAD6",
X"BADF2F",
X"BBF552",
X"BD0D38",
X"BE26D9",
X"BF422E",
X"C05F30",
X"C17DD8",
X"C29E1E",
X"C3BFFA",
X"C4E365",
X"C60858",
X"C72ECA",
X"C856B5",
X"C98011",
X"CAAAD6",
X"CBD6FB",
X"CD047B",
X"CE334C",
X"CF6367",
X"D094C3",
X"D1C75A",
X"D2FB23",
X"D43016",
X"D5662C",
X"D69D5B",
X"D7D59D",
X"D90EE9",
X"DA4936",
X"DB847E",
X"DCC0B7",
X"DDFDD9",
X"DF3BDD",
X"E07ABA",
X"E1BA67",
X"E2FADD",
X"E43C13",
X"E57E01",
X"E6C09F",
X"E803E4",
X"E947C8",
X"EA8C42",
X"EBD14A",
X"ED16D8",
X"EE5CE4",
X"EFA364",
X"F0EA50",
X"F231A1",
X"F3794C",
X"F4C14B",
X"F60995",
X"F75220",
X"F89AE4",
X"F9E3DA",
X"FB2CF8",
X"FC7636",
X"FDBF8C",
X"FF08F0",
X"00525A",
X"019BC3",
X"02E521",
X"042E6C",
X"05779B",
X"06C0A6",
X"080985",
X"09522E",
X"0A9A99",
X"0BE2BE",
X"0D2A94",
X"0E7213",
X"0FB933",
X"10FFEA",
X"124631",
X"138BFF",
X"14D14B",
X"16160D",
X"175A3D",
X"189DD3",
X"19E0C5",
X"1B230C",
X"1C649F",
X"1DA576",
X"1EE589",
X"2024CF",
X"216341",
X"22A0D5",
X"23DD84",
X"251945",
X"265410",
X"278DDE",
X"28C6A6",
X"29FE5F",
X"2B3503",
X"2C6A88",
X"2D9EE7",
X"2ED218",
X"300413",
X"3134D0",
X"326447",
X"339270",
X"34BF43",
X"35EAB9",
X"3714CA",
X"383D6F",
X"39649F",
X"3A8A52",
X"3BAE82",
X"3CD127",
X"3DF239",
X"3F11B0",
X"402F86",
X"414BB2",
X"42662F",
X"437EF3",
X"4495F8",
X"45AB38",
X"46BEA9",
X"47D046",
X"48E008",
X"49EDE7",
X"4AF9DC",
X"4C03E0",
X"4D0BED",
X"4E11FC",
X"4F1606",
X"501803",
X"5117EF",
X"5215C1",
X"531174",
X"540B00",
X"550260",
X"55F78C",
X"56EA80",
X"57DB33",
X"58C9A1",
X"59B5C3",
X"5A9F92",
X"5B870A",
X"5C6C23",
X"5D4ED8",
X"5E2F22",
X"5F0CFE",
X"5FE863",
X"60C14D",
X"6197B7",
X"626B9A",
X"633CF1",
X"640BB7",
X"64D7E6",
X"65A17A",
X"66686C",
X"672CB8",
X"67EE58",
X"68AD49",
X"696984",
X"6A2304",
X"6AD9C6",
X"6B8DC4",
X"6C3EFA",
X"6CED63",
X"6D98FA",
X"6E41BB",
X"6EE7A2",
X"6F8AAB",
X"702AD1",
X"70C810",
X"716263",
X"71F9C8",
X"728E3A",
X"731FB6",
X"73AE36",
X"7439B9",
X"74C23A",
X"7547B5",
X"75CA28",
X"76498E",
X"76C5E5",
X"773F2A",
X"77B558",
X"78286E",
X"789868",
X"790543",
X"796EFC",
X"79D592",
X"7A3900",
X"7A9945",
X"7AF65D",
X"7B5048",
X"7BA701",
X"7BFA88",
X"7C4AD9",
X"7C97F4",
X"7CE1D5",
X"7D287B",
X"7D6BE3",
X"7DAC0E",
X"7DE8F7",
X"7E229F",
X"7E5904",
X"7E8C23",
X"7EBBFD",
X"7EE88F",
X"7F11D8",
X"7F37D8",
X"7F5A8E",
X"7F79F7",
X"7F9615",
X"7FAEE5",
X"7FC468",
X"7FD69C",
X"7FE582",
X"7FF119",
X"7FF960",
X"7FFE58");
begin
	cosx <= cosxrom(address);
end cos625_24bit_ARCH;



