library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity sin625_24bit is
	port( address : IN INTEGER := 0;
		 sinx : OUT std_logic_vector (23 downto 0));
end sin625_24bit;

architecture sin625_24bit_ARCH of sin625_24bit is
	type sinromarray is array (0 to 624) of std_logic_vector (23 downto 0);
	constant sinxrom : sinromarray := (
X"000000",
X"01496A",
X"0292CB",
X"03DC1C",
X"052553",
X"066E67",
X"07B752",
X"090009",
X"0A4884",
X"0B90BC",
X"0CD8A7",
X"0E203C",
X"0F6775",
X"10AE47",
X"11F4AA",
X"133A97",
X"148004",
X"15C4EA",
X"17093F",
X"184CFC",
X"199018",
X"1AD28B",
X"1C144C",
X"1D5553",
X"1E9597",
X"1FD511",
X"2113B9",
X"225185",
X"238E6E",
X"24CA6B",
X"260575",
X"273F83",
X"28788D",
X"29B08B",
X"2AE774",
X"2C1D42",
X"2D51EB",
X"2E8569",
X"2FB7B2",
X"30E8BF",
X"321888",
X"334705",
X"34742F",
X"359FFD",
X"36CA68",
X"37F368",
X"391AF6",
X"3A4109",
X"3B659B",
X"3C88A3",
X"3DAA1A",
X"3EC9F9",
X"3FE838",
X"4104D0",
X"421FB9",
X"4338EC",
X"445061",
X"456613",
X"4679F8",
X"478C0B",
X"489C44",
X"49AA9C",
X"4AB70D",
X"4BC18E",
X"4CCA19",
X"4DD0A8",
X"4ED534",
X"4FD7B5",
X"50D826",
X"51D67F",
X"52D2BA",
X"53CCD1",
X"54C4BC",
X"55BA76",
X"56ADF9",
X"579F3D",
X"588E3D",
X"597AF2",
X"5A6556",
X"5B4D64",
X"5C3316",
X"5D1664",
X"5DF74A",
X"5ED5C2",
X"5FB1C5",
X"608B4F",
X"616259",
X"6236DE",
X"6308D9",
X"63D843",
X"64A519",
X"656F54",
X"6636EF",
X"66FBE5",
X"67BE31",
X"687DCD",
X"693AB6",
X"69F4E6",
X"6AAC58",
X"6B6107",
X"6C12EF",
X"6CC20C",
X"6D6E58",
X"6E17CF",
X"6EBE6D",
X"6F622E",
X"70030D",
X"70A106",
X"713C15",
X"71D436",
X"726965",
X"72FB9E",
X"738ADE",
X"741720",
X"74A062",
X"75269F",
X"75A9D4",
X"7629FE",
X"76A719",
X"772122",
X"779817",
X"780BF3",
X"787CB4",
X"78EA57",
X"7954D9",
X"79BC38",
X"7A2070",
X"7A817F",
X"7ADF63",
X"7B3A1A",
X"7B91A0",
X"7BE5F3",
X"7C3712",
X"7C84FA",
X"7CCFAA",
X"7D171F",
X"7D5B57",
X"7D9C51",
X"7DDA0B",
X"7E1484",
X"7E4BB9",
X"7E7FAA",
X"7EB055",
X"7EDDB9",
X"7F07D5",
X"7F2EA7",
X"7F522F",
X"7F726C",
X"7F8F5D",
X"7FA900",
X"7FBF56",
X"7FD25F",
X"7FE218",
X"7FEE82",
X"7FF79E",
X"7FFD69",
X"7FFFE5",
X"7FFF11",
X"7FFAED",
X"7FF37A",
X"7FE8B7",
X"7FDAA5",
X"7FC944",
X"7FB495",
X"7F9C98",
X"7F814E",
X"7F62B7",
X"7F40D5",
X"7F1BA7",
X"7EF330",
X"7EC770",
X"7E9868",
X"7E661A",
X"7E3087",
X"7DF7B0",
X"7DBB96",
X"7D7C3C",
X"7D39A3",
X"7CF3CC",
X"7CAAB9",
X"7C5E6D",
X"7C0EE9",
X"7BBC30",
X"7B6643",
X"7B0D24",
X"7AB0D7",
X"7A515D",
X"79EEB9",
X"7988ED",
X"791FFC",
X"78B3E9",
X"7844B7",
X"77D268",
X"775CFF",
X"76E480",
X"7668EE",
X"75EA4B",
X"75689B",
X"74E3E1",
X"745C21",
X"73D15F",
X"73439D",
X"72B2E0",
X"721F2C",
X"718883",
X"70EEEB",
X"705266",
X"6FB2FA",
X"6F10AA",
X"6E6B7A",
X"6DC36E",
X"6D188C",
X"6C6AD7",
X"6BBA55",
X"6B0708",
X"6A50F7",
X"699825",
X"68DC99",
X"681E55",
X"675D60",
X"6699BF",
X"65D376",
X"650A8A",
X"643F01",
X"6370E0",
X"62A02D",
X"61CCEC",
X"60F724",
X"601ED9",
X"5F4412",
X"5E66D4",
X"5D8724",
X"5CA509",
X"5BC089",
X"5AD9A9",
X"59F06F",
X"5904E1",
X"581706",
X"5726E3",
X"56347F",
X"553FE0",
X"54490C",
X"53500B",
X"5254E1",
X"515796",
X"505830",
X"4F56B6",
X"4E532F",
X"4D4DA1",
X"4C4613",
X"4B3C8C",
X"4A3112",
X"4923AD",
X"481464",
X"47033D",
X"45F03F",
X"44DB73",
X"43C4DF",
X"42AC89",
X"41927A",
X"4076B9",
X"3F594D",
X"3E3A3D",
X"3D1991",
X"3BF751",
X"3AD383",
X"39AE2F",
X"38875E",
X"375F16",
X"36355F",
X"350A42",
X"33DDC5",
X"32AFF0",
X"3180CC",
X"305060",
X"2F1EB4",
X"2DEBD0",
X"2CB7BC",
X"2B827F",
X"2A4C22",
X"2914AE",
X"27DC29",
X"26A29C",
X"25680F",
X"242C8A",
X"22F016",
X"21B2BB",
X"207480",
X"1F356E",
X"1DF58E",
X"1CB4E7",
X"1B7382",
X"1A3167",
X"18EE9F",
X"17AB32",
X"166727",
X"152289",
X"13DD5E",
X"1297B0",
X"115187",
X"100AEB",
X"0EC3E5",
X"0D7C7D",
X"0C34BB",
X"0AECA9",
X"09A44F",
X"085BB4",
X"0712E2",
X"05C9E2",
X"0480BB",
X"033776",
X"01EE1C",
X"00A4B5",
X"FF5B4B",
X"FE11E4",
X"FCC88A",
X"FB7F45",
X"FA361E",
X"F8ED1E",
X"F7A44C",
X"F65BB1",
X"F51357",
X"F3CB45",
X"F28383",
X"F13C1B",
X"EFF515",
X"EEAE79",
X"ED6850",
X"EC22A2",
X"EADD77",
X"E998D9",
X"E854CE",
X"E71161",
X"E5CE99",
X"E48C7E",
X"E34B19",
X"E20A72",
X"E0CA92",
X"DF8B80",
X"DE4D45",
X"DD0FEA",
X"DBD376",
X"DA97F1",
X"D95D64",
X"D823D7",
X"D6EB52",
X"D5B3DE",
X"D47D81",
X"D34844",
X"D21430",
X"D0E14C",
X"CFAFA0",
X"CE7F34",
X"CD5010",
X"CC223B",
X"CAF5BE",
X"C9CAA1",
X"C8A0EA",
X"C778A2",
X"C651D1",
X"C52C7D",
X"C408AF",
X"C2E66F",
X"C1C5C3",
X"C0A6B3",
X"BF8947",
X"BE6D86",
X"BD5377",
X"BC3B21",
X"BB248D",
X"BA0FC1",
X"B8FCC3",
X"B7EB9C",
X"B6DC53",
X"B5CEEE",
X"B4C374",
X"B3B9ED",
X"B2B25F",
X"B1ACD1",
X"B0A94A",
X"AFA7D0",
X"AEA86A",
X"ADAB1F",
X"ACAFF5",
X"ABB6F4",
X"AAC020",
X"A9CB81",
X"A8D91D",
X"A7E8FA",
X"A6FB1F",
X"A60F91",
X"A52657",
X"A43F77",
X"A35AF7",
X"A278DC",
X"A1992C",
X"A0BBEE",
X"9FE127",
X"9F08DC",
X"9E3314",
X"9D5FD3",
X"9C8F20",
X"9BC0FF",
X"9AF576",
X"9A2C8A",
X"996641",
X"98A2A0",
X"97E1AB",
X"972367",
X"9667DB",
X"95AF09",
X"94F8F8",
X"9445AB",
X"939529",
X"92E774",
X"923C92",
X"919486",
X"90EF56",
X"904D06",
X"8FAD9A",
X"8F1115",
X"8E777D",
X"8DE0D4",
X"8D4D20",
X"8CBC63",
X"8C2EA1",
X"8BA3DF",
X"8B1C1F",
X"8A9765",
X"8A15B5",
X"899712",
X"891B80",
X"88A301",
X"882D98",
X"87BB49",
X"874C17",
X"86E004",
X"867713",
X"861147",
X"85AEA3",
X"854F29",
X"84F2DC",
X"8499BD",
X"8443D0",
X"83F117",
X"83A193",
X"835547",
X"830C34",
X"82C65D",
X"8283C4",
X"82446A",
X"820850",
X"81CF79",
X"8199E6",
X"816798",
X"813890",
X"810CD0",
X"80E459",
X"80BF2B",
X"809D49",
X"807EB2",
X"806368",
X"804B6B",
X"8036BC",
X"80255B",
X"801749",
X"800C86",
X"800513",
X"8000EF",
X"80001B",
X"800297",
X"800862",
X"80117E",
X"801DE8",
X"802DA1",
X"8040AA",
X"805700",
X"8070A3",
X"808D94",
X"80ADD1",
X"80D159",
X"80F82B",
X"812247",
X"814FAB",
X"818056",
X"81B447",
X"81EB7C",
X"8225F5",
X"8263AF",
X"82A4A9",
X"82E8E1",
X"833056",
X"837B06",
X"83C8EE",
X"841A0D",
X"846E60",
X"84C5E6",
X"85209D",
X"857E81",
X"85DF90",
X"8643C8",
X"86AB27",
X"8715A9",
X"87834C",
X"87F40D",
X"8867E9",
X"88DEDE",
X"8958E7",
X"89D602",
X"8A562C",
X"8AD961",
X"8B5F9E",
X"8BE8E0",
X"8C7522",
X"8D0462",
X"8D969B",
X"8E2BCA",
X"8EC3EB",
X"8F5EFA",
X"8FFCF3",
X"909DD2",
X"914193",
X"91E831",
X"9291A8",
X"933DF4",
X"93ED11",
X"949EF9",
X"9553A8",
X"960B1A",
X"96C54A",
X"978233",
X"9841CF",
X"99041B",
X"99C911",
X"9A90AC",
X"9B5AE7",
X"9C27BD",
X"9CF727",
X"9DC922",
X"9E9DA7",
X"9F74B1",
X"A04E3B",
X"A12A3E",
X"A208B6",
X"A2E99C",
X"A3CCEA",
X"A4B29C",
X"A59AAA",
X"A6850E",
X"A771C3",
X"A860C3",
X"A95207",
X"AA458A",
X"AB3B44",
X"AC332F",
X"AD2D46",
X"AE2981",
X"AF27DA",
X"B0284B",
X"B12ACC",
X"B22F58",
X"B335E7",
X"B43E72",
X"B548F3",
X"B65564",
X"B763BC",
X"B873F5",
X"B98608",
X"BA99ED",
X"BBAF9F",
X"BCC714",
X"BDE047",
X"BEFB30",
X"C017C8",
X"C13607",
X"C255E6",
X"C3775D",
X"C49A65",
X"C5BEF7",
X"C6E50A",
X"C80C98",
X"C93598",
X"CA6003",
X"CB8BD1",
X"CCB8FB",
X"CDE778",
X"CF1741",
X"D0484E",
X"D17A97",
X"D2AE15",
X"D3E2BE",
X"D5188C",
X"D64F75",
X"D78773",
X"D8C07D",
X"D9FA8B",
X"DB3595",
X"DC7192",
X"DDAE7B",
X"DEEC47",
X"E02AEF",
X"E16A69",
X"E2AAAD",
X"E3EBB4",
X"E52D75",
X"E66FE8",
X"E7B304",
X"E8F6C1",
X"EA3B16",
X"EB7FFC",
X"ECC569",
X"EE0B56",
X"EF51B9",
X"F0988B",
X"F1DFC4",
X"F32759",
X"F46F44",
X"F5B77C",
X"F6FFF7",
X"F848AE",
X"F99199",
X"FADAAD",
X"FC23E4",
X"FD6D35",
X"FEB696");
begin
	sinx <= sinxrom(address);
end sin625_24bit_ARCH;


